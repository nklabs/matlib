// Square root step

// Copyright 2023 NK Labs, LLC

// Permission is hereby granted, free of charge, to any person obtaining a
// copy of this software and associated documentation files (the
// "Software"), to deal in the Software without restriction, including
// without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to permit
// persons to whom the Software is furnished to do so, subject to the
// following conditions:

// The above copyright notice and this permission notice shall be included
// in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
// OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. 
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY
// CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT
// OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR
// THE USE OR OTHER DEALINGS IN THE SOFTWARE.

module sqrt_step
  (
  fixedp g, // Fixed point parameters and common ports

  input [g.WIDTH:0] r_in,
  input [g.WIDTH:0] b_in,
  input [g.WIDTH:0] q_in,

  output reg [g.WIDTH:0] r,
  output reg [g.WIDTH:0] b,
  output reg [g.WIDTH:0] q
  );

wire [g.WIDTH:0] newr = r_in - (q_in + b_in);

always @(posedge g.clk)
  begin
    if (r_in >= q_in + b_in)
      begin
        r <= { newr[g.WIDTH-1:0], 1'd0 };
        q <= q_in + { b_in[g.WIDTH-1:0], 1'd0 };
      end
    else
      begin
        r <= { r_in[g.WIDTH-1:0], 1'd0 };
        q <= q_in;
      end
    b <= { 1'd0, b_in[g.WIDTH:1] };
  end

endmodule
