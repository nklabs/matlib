// Return element of vector with maximum absolute value

// Copyright 2023 NK Labs, LLC

// Permission is hereby granted, free of charge, to any person obtaining a
// copy of this software and associated documentation files (the
// "Software"), to deal in the Software without restriction, including
// without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to permit
// persons to whom the Software is furnished to do so, subject to the
// following conditions:

// The above copyright notice and this permission notice shall be included
// in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
// OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. 
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY
// CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT
// OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR
// THE USE OR OTHER DEALINGS IN THE SOFTWARE.

module vecmaxmag
 #(
  parameter COLS = 1
) (
  fixedp g, // Fixed point parameters and common ports

  input signed [COLS:1][g.WIDTH-1:0] a,
  output logic [g.WIDTH-1:0] f
  );

logic signed [g.WIDTH-1:0] themax;
logic signed [g.WIDTH-1:0] absthemax;
logic signed [g.WIDTH-1:0] tmp;

always @(posedge g.clk)
  begin
    f <= themax;
  end

always @*
  begin
    themax = a[1];
    if (a[1][g.WIDTH-1])
      absthemax = -a[1];
    else
      absthemax = a[1];

    for (int i = 2; i <= COLS; i = i + 1)
      begin
        if (a[i][g.WIDTH-1])
          tmp = -a[i];
        else
          tmp = a[i];
        if (tmp > absthemax)
          begin
            absthemax = tmp;
            themax = a[i];
          end
      end
  end

endmodule
